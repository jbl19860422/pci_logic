LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY DIV IS
PORT
(
	RST		:IN STD_LOGIC;
	INCLK0	:IN	STD_LOGIC;	--����ʱ��
	OUTCLK0	:INOUT	STD_LOGIC;--����Ƶ
	OUTCLK1	:INOUT	STD_LOGIC;--�ķ�Ƶ
	OUTCLK2	:INOUT	STD_LOGIC--�˷�Ƶ
);
END DIV;

ARCHITECTURE STR OF DIV IS

BEGIN

PROCESS (RST,INCLK0)
BEGIN
	IF(RST = '0') THEN
		OUTCLK0 <= '0';
	ELSIF(INCLK0'EVENT AND INCLK0 = '1') THEN
			OUTCLK0 <= NOT OUTCLK0;
	END IF;
END PROCESS;

PROCESS(RST,OUTCLK0)
BEGIN
	IF(RST = '0') THEN
		OUTCLK1 <= '0';
	ELSIF(OUTCLK0'EVENT AND OUTCLK0 = '1') THEN
			OUTCLK1 <= NOT OUTCLK1;
	END IF;
END PROCESS;

PROCESS(RST,OUTCLK1)
BEGIN
	IF(RST = '0') THEN
		OUTCLK2 <= '0';
	ELSIF(OUTCLK1'EVENT AND OUTCLK1 = '1') THEN
			OUTCLK2 <= NOT OUTCLK2;
	END IF;
END PROCESS;

END STR;