LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
PACKAGE Type_Pkg IS
TYPE Array_Addr4 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(3 DOWNTO 0);
TYPE Array_Addr5 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(4 DOWNTO 0);
TYPE Array_Channel IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(4 DOWNTO 0);
TYPE A_V37 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(36 DOWNTO 0);
TYPE A_V6 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(5 DOWNTO 0);
TYPE A_V32 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
TYPE A_V20 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(19 DOWNTO 0);
TYPE A_V28 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(27 DOWNTO 0);
TYPE A_V54 IS ARRAY(NATURAL RANGE<>) OF STD_LOGIC_VECTOR(53 DOWNTO 0);
END Type_Pkg;