LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;


ENTITY DIV_2 IS
PORT
(
	RST		:IN STD_LOGIC;
	En			:IN STD_LOGIC;
	INCLK0	:IN STD_LOGIC;	--����ʱ��
	OUTCLK0	:OUT	STD_LOGIC
);
END DIV_2;

ARCHITECTURE STR OF DIV_2 IS
SIGNAL OUTCLK0_Tmp:STD_LOGIC;
BEGIN

PROCESS (RST,En, INCLK0)
BEGIN
	IF(RST = '0') OR En = '0' THEN
		OUTCLK0_Tmp <= '0';
	ELSIF(INCLK0'EVENT AND INCLK0 = '1') THEN
		IF En = '1' THEN
			OUTCLK0_Tmp <= NOT OUTCLK0_Tmp;
		ELSE
			OUTCLK0_Tmp <= '0';
		END IF;
	END IF;
END PROCESS;
OUTCLK0 <= OUTCLK0_Tmp;
END STR;