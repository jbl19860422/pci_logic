PLL_80_inst : PLL_80 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
