LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE DEFINE IS
--	TYPE STATUSSET IS (IDLE_NOR,BUSY,SDATA,TURNAROUND);
	
	CONSTANT IO            : STD_LOGIC := '1';
	CONSTANT MEM           : STD_LOGIC := '0'; 
	CONSTANT IOMEM         : STD_LOGIC_VECTOR(5 DOWNTO 0) := "00000" & IO;

	CONSTANT Device_ID     : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"0001"; 
	CONSTANT Vendor_ID     : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"1103";
	CONSTANT CFCSTATUS     : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"0400";	  -- Slow Devsel
	CONSTANT CFGCOMMAND    : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"0001";    -- IO Access
	CONSTANT Class_Code    : STD_LOGIC_VECTOR(23 DOWNTO 0) := X"028000";  -- Network Controller
    CONSTANT Revision_ID   : STD_LOGIC_VECTOR(7  DOWNTO 0) := X"01";		
	CONSTANT BIST          : STD_LOGIC_VECTOR(7  DOWNTO 0) := X"00";      -- Not Support BIST
	CONSTANT Header_Type   : STD_LOGIC_VECTOR(7  DOWNTO 0) := X"00";
	CONSTANT Latency_Timer : STD_LOGIC_VECTOR(7  DOWNTO 0) := X"00";      -- Not Support in Slave
	CONSTANT Cache_Size    : STD_LOGIC_VECTOR(7  DOWNTO 0) := X"00";	  -- Not Cache Access
	CONSTANT Int_Pin       : STD_LOGIC_VECTOR(7  DOWNTO 0) := X"01";      -- Use INTA
	
	CONSTANT NULL8         : STD_LOGIC_VECTOR(7  DOWNTO 0) := X"00";
	CONSTANT NULL16        : STD_LOGIC_VECTOR(15 DOWNTO 0) := X"0000";
	CONSTANT NULL24        : STD_LOGIC_VECTOR(23 DOWNTO 0) := X"000000";
	CONSTANT NULL32        : STD_LOGIC_VECTOR(31 DOWNTO 0) := X"00000000";
	
	CONSTANT High8         : STD_LOGIC_VECTOR(7  DOWNTO 0) := "ZZZZZZZZ";
	CONSTANT High16        : STD_LOGIC_VECTOR(15 DOWNTO 0) := "ZZZZZZZZZZZZZZZZ";
	CONSTANT High24        : STD_LOGIC_VECTOR(23 DOWNTO 0) := "ZZZZZZZZZZZZZZZZZZZZZZZZ";
	CONSTANT High32        : STD_LOGIC_VECTOR(31 DOWNTO 0) := "ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ";

END DEFINE;

PACKAGE BODY DEFINE IS
END DEFINE;